/nfs/site/disks/vmisd_vclp_efficiency/rcg/test/cadence/rcgFlow/AsicMethadology/riscvCoreSyntaCore1/ramInputs/sram_32_1024.lef