/home/cadence/Documents/raksha/AsicMethadology/technology/45/lef/MEM2_128X32.lef