/nfs/site/disks/vmisd_vclp_efficiency/rcg/test/cadence/rcgFlow/AsicMethadology/riscvCoreSyntaCore1/ramInputs/scr1_pipe_top.lef