/home/cadence/Documents/raksha/AsicMethadology/technology/45/lef/MEM1_256X32.lef