/nfs/site/disks/vmisd_vclp_efficiency/rcg/test/cadence/venvRcg/AsicMethadology/riscvCoreSyntaCore1/ramInputs/i2c_top.lef