/home/cadence/Documents/raksha/AsicMethadology/technology/45/lef/pads.lef