/nfs/site/disks/vmisd_vclp_efficiency/rcg/test/cadence/rcgFlow/AsicMethadology/technology/45/lef/pdkIO.lef