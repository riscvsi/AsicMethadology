/home/cadence/Documents/raksha/AsicMethadology/technology/45/lef/gsclib045.fixed2.lef